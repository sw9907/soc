module adder(
		input			a,
		input 			b,
		output wire 	y
		);

assign y = a + b;

endmodule
